/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_teletext.cdl
 * @brief Testbench for teletext decoder module
 *
 * This is a simple testbench for the teletext decoder.
 */
/*a Includes */
include "apb::csr.h"
include "bbc_types.h"
include "bbc_submodules.h"

/*a Module */
module tb_bbc_with_shm_display( clock system_clk,
                                clock system_clk_div_2,
                                clock video_clk,
                                input bit reset_n
)
{

    /*b Nets */
    default clock system_clk;
    default reset active_low reset_n;
    net t_csr_request csr_request;
    net t_csr_response csr_response;
    net t_bbc_micro_sram_request   host_sram_request;
    net t_bbc_micro_sram_response host_sram_response;
    net t_bbc_display_sram_write display_sram_write;
    instances : {
        bbc_micro_with_rams bbc( clk<-system_clk,
                       video_clk<-video_clk,

                       reset_n <= reset_n,
                       host_sram_request <= host_sram_request,
                       csr_request <= csr_request,
                       display_sram_write => display_sram_write,
                       host_sram_response => host_sram_response,
                       csr_response => csr_response );
        bbc_display display( clk <- system_clk_div_2,
                             host_sram_request => host_sram_request,
                             csr_request => csr_request,
                             display_sram_write <= display_sram_write,
                             host_sram_response <= host_sram_response,
                             csr_response <= csr_response );
    }
}

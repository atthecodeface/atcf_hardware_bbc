/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file   bbc_micro_de1_cl_bbc.cdl
 * @brief  BBC microcomputer with RAMs for the CL DE1 + daughterboard
 *
 * CDL module containing the BBC microcomputer with RAMs and associated logic
 * for the Cambridge University Computer Laboratory DE1 + daughterboard system.
 *
 */
/*a Includes */
include "bbc::bbc_types.h"
include "bbc::bbc_submodules.h"
include "std::srams.h"
include "video::framebuffer_modules.h"

/*a Module */
module bbc_micro_de1_cl_bbc( clock clk          "50MHz clock from DE1 clock generator",
                             clock video_clk    "9MHz clock from PLL, derived from 50MHz",
                             input bit reset_n  "hard reset from a pin - a key on DE1",
                             input bit bbc_reset_n,
                             input bit framebuffer_reset_n,
                             output t_bbc_clock_control clock_control,
                             input t_bbc_keyboard bbc_keyboard,
                             output t_video_bus video_bus,
                             input t_csr_request csr_request,
                             output t_csr_response csr_response
    )
{

    net t_bbc_display display;
    net t_bbc_floppy_op floppy_op;
    net  t_bbc_floppy_response floppy_response;

    net t_bbc_clock_status clock_status;
    net t_bbc_clock_control clock_control;

    clocked clock clk reset active_low reset_n t_csr_response csr_response={*=0};
    comb t_csr_response combined_csr_response;
    net t_csr_response clocking_csr_response;
    net t_csr_response display_sram_csr_response;
    net t_csr_response floppy_sram_csr_response;
    net t_csr_response framebuffer_csr_response;
    net t_video_bus video_bus;

    net t_bbc_floppy_sram_request floppy_sram_request;
    net t_bbc_display_sram_write display_sram_write;

    comb t_bbc_micro_sram_request  bbc_micro_host_sram_request;
    net  t_bbc_micro_sram_response bbc_micro_host_sram_response;
    
    gated_clock clock clk active_high enable_clk_2MHz_video   clk_2MHz_video_clock "Clock that mirrors 2MHz falling -  video data from RAM is valid at this edge, so used by CRTC, SAA5050 latches, SAA5050, vidproc";
    gated_clock clock clk active_high enable_cpu_clk          clk_cpu  "6502 clock, >=2MHz but extended when accessing 1MHz peripherals";
    comb bit enable_clk_2MHz_video;
    comb bit enable_cpu_clk;

    net bit[32] floppy_sram_read_data;
    clocked clock clk_cpu reset active_low reset_n bit floppy_sram_reading=0;
    clocked clock clk_cpu reset active_low reset_n t_bbc_floppy_sram_request floppy_sram_request_r={*=0};
    clocked clock clk_cpu reset active_low reset_n t_bbc_floppy_sram_response floppy_sram_response={*=0};

    /*b BBC Micro instantiations */
    bbc_micro_instantiations: {
        bbc_micro_host_sram_request = {*=0};
        enable_cpu_clk        = clock_control.enable_cpu;
        enable_clk_2MHz_video = clock_control.enable_2MHz_video;
        combined_csr_response  = clocking_csr_response;
        combined_csr_response |= display_sram_csr_response;
        combined_csr_response |= floppy_sram_csr_response;
        combined_csr_response |= framebuffer_csr_response;
        csr_response <= combined_csr_response;
        bbc_micro_clocking clocking( clk <- clk,
                                     reset_n <= reset_n,
                                     clock_status <= clock_status,
                                     clock_control => clock_control,
                                     csr_request <= csr_request,
                                     csr_response => clocking_csr_response );

        bbc_micro bbc(clk <- clk,
                      reset_n <= bbc_reset_n,
                      clock_control <= clock_control,
                      clock_status  => clock_status,
                      keyboard <= bbc_keyboard,
                      display => display,
                      floppy_op => floppy_op,
                      floppy_response <= floppy_response,
                      host_sram_request <= bbc_micro_host_sram_request,
                      host_sram_response => bbc_micro_host_sram_response
            );
    
        bbc_display_sram display_sram( clk <- clk_2MHz_video_clock,
                                       reset_n <= reset_n,
                                       display <= display,
                                       sram_write => display_sram_write,
                                       csr_request <= csr_request,
                                       csr_response => display_sram_csr_response
            );

        bbc_floppy_sram floppy_sram( clk <- clk_cpu, // FDC interacts with floppy at cpu clock
                                     reset_n <= reset_n,
                                     floppy_op <= floppy_op,
                                     csr_request <= csr_request,
                                     floppy_response => floppy_response,
                                     sram_request => floppy_sram_request,
                                     sram_response <= floppy_sram_response,
                                     csr_response => floppy_sram_csr_response
            );

    }

    /*b SRAMs for floppy and framebuffers */
    comb t_sram_access_req display_sram_access_req;
    floppy_and_framebuffer: {
        se_sram_srw_32768x32 floppy(sram_clock <- clk_cpu,
                                    select         <= floppy_sram_request_r.enable && !floppy_sram_reading,
                                    read_not_write <= floppy_sram_request_r.read_not_write,
                                    write_enable   <= !floppy_sram_request_r.read_not_write,
                                    address        <= floppy_sram_request_r.address[15;0],
                                    write_data     <= floppy_sram_request_r.write_data[32;0],
                                    data_out       => floppy_sram_read_data );
        floppy_sram_request_r    <= floppy_sram_request;
        floppy_sram_reading      <= (floppy_sram_request_r.enable && !floppy_sram_reading) && floppy_sram_request_r.read_not_write;
        floppy_sram_response.ack  <= floppy_sram_request.enable;
        floppy_sram_response.read_data_valid <= floppy_sram_reading;
        floppy_sram_response.read_data       <= floppy_sram_read_data;

        display_sram_access_req = {*=0};
        display_sram_access_req.valid      = display_sram_write.enable;
        display_sram_access_req.address    = bundle(16b0,display_sram_write.address);
        display_sram_access_req.write_data = bundle(16b0,display_sram_write.data);
        framebuffer fb( csr_clk <- clk_cpu,
                        sram_clk <- clk_2MHz_video_clock,
                        video_clk <- video_clk,
                        reset_n <= framebuffer_reset_n,
                        video_bus => video_bus,
                        display_sram_write <= display_sram_access_req,
                        csr_request <= csr_request,
                        csr_response => framebuffer_csr_response
            );
                        
    }

    /*b All done */
}
